carrt